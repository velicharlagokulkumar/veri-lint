module counter #( 
    parameter WIDTH = 8
)(
    input clk, 
    input reset,
    output logic [WIDTH-1 : 0] out
);

  always @(posedge clk) begin
    if (reset)
      out <= 0;
    else
      out <= out + 1;
    end

endmodule