module test();
    initial begin
        $display("Hello, SystemVerilog!");
    end
endmodule
