module tb;
    test uut();
    initial begin
        #10;
        $finish;
    end
endmodule
